module main (
	
	);

endmodule
